//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4_2
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//                                          
// DESCRIPTION: This test extends test_top and makes 
//    changes to test_top using the UVM factory type_override:
//
//    Test scenario: 
//      This is a template test that can be used to create future tests.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

class singleADDinstr_test extends test_top;

  `uvm_component_utils( singleADDinstr_test );

  function new( string name = "", uvm_component parent = null );
    super.new( name, parent );
  endfunction

  virtual function void build_phase(uvm_phase phase);
    // The factory override below replaces the lc3_bench_sequence_base 
    // sequence with the register_test_sequence.
    //lc3_bench_sequence_base::type_id::set_type_override(register_test_sequence::get_type());

    //Harry: debug message
    `uvm_info("singleADDinstr_test", "Harry-> imem_responder_singleADDinstr_sequence overridding imem_responder_sequence(base)...", UVM_HIGH)

    //Harry: Override the instruction memory responder with our single ADD instruction program
    set_type_override_by_type(
      imem_responder_sequence::get_type(),
      imem_responder_singleADDinstr_sequence::get_type()
    );
    // Execute the build_phase of test_top AFTER all factory overrides have been created.
    super.build_phase(phase);
  endfunction

  virtual task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    `uvm_info("SINGLEADDINSTR_TEST", "===== LC3 SINGLE ADD INSTRUCTION TEST START =====", UVM_LOW)
    super.run_phase(phase); // let uvmf_test_base start LC3_bench_sequence_base
    #1us; //Harry->question: how long should we run the simulation?
    `uvm_info("SINGLEADDINSTR_TEST", "===== LC3 SINGLE ADD INSTRUCTION TEST COMPLETE =====", UVM_LOW)
    phase.drop_objection(this);
  endtask

  virtual function void end_of_elaboration_phase(uvm_phase phase);
    super.end_of_elaboration_phase(phase);
    // pragma uvmf custom register_test_scoreboard_control begin

    // These UVMF scoreboards may need to be disabled for the register test.  
    
    // environment.fetch_env.fetch_scoreboard.disable_scoreboard();
    // environment.fetch_env.fetch_scoreboard.disable_end_of_test_activity_check();
    
    // environment.decode_env.decode_scoreboard.disable_scoreboard();
    // environment.decode_env.decode_scoreboard.disable_end_of_test_activity_check();
    
    // environment.execute_env.execute_scoreboard.disable_scoreboard();
    // environment.execute_env.execute_scoreboard.disable_end_of_test_activity_check();
    
    // environment.writeback_env.writeback_scoreboard.disable_scoreboard();
    // environment.writeback_env.writeback_scoreboard.disable_end_of_test_activity_check();
    
    // environment.memaccess_env.memaccess_scoreboard.disable_scoreboard();
    // environment.memaccess_env.memaccess_scoreboard.disable_end_of_test_activity_check();
    
    // environment.controller_env.controller_scoreboard.disable_scoreboard();
    // environment.controller_env.controller_scoreboard.disable_end_of_test_activity_check();
    
    // pragma uvmf custom register_test_scoreboard_control end
  endfunction

endclass

// pragma uvmf custom external begin
// pragma uvmf custom external end

