module  hvl_qvip_agents 
      #(
        string HDL_BFM_SCOPE = "",
        string HVL_AGENT_SCOPE = ""
       );

  initial begin
    $display("Hello World from QVIP hvl");
  end

endmodule

