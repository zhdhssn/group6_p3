//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4_2
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//
//----------------------------------------------------------------------
//
// DESCRIPTION: This analysis component contains analysis_exports for receiving
//   data and analysis_ports for sending data.
// 
//   This analysis component has the following analysis_exports that receive the 
//   listed transaction type.
//   
//   decode_in_ae receives transactions of type  decode_in_transaction
//
//   This analysis component has the following analysis_ports that can broadcast 
//   the listed transaction type.
//
//  decode_out_ap broadcasts transactions of type decode_out_transaction
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
import lc3_prediction_pkg::*;

class decode_predictor #(
  type CONFIG_T,
  type BASE_T = uvm_component
  )
 extends BASE_T;

  // Factory registration of this class
  `uvm_component_param_utils( decode_predictor #(
                              CONFIG_T,
                              BASE_T
                              )
)


  // Instantiate a handle to the configuration of the environment in which this component resides
  CONFIG_T configuration;

  
  // Instantiate the analysis exports
  uvm_analysis_imp_decode_in_ae #(decode_in_transaction, decode_predictor #(
                              .CONFIG_T(CONFIG_T),
                              .BASE_T(BASE_T)
                              )
) decode_in_ae;

  
  // Instantiate the analysis ports
  uvm_analysis_port #(decode_out_transaction) decode_out_ap;


  // Transaction variable for predicted values to be sent out decode_out_ap
  // Once a transaction is sent through an analysis_port, another transaction should
  // be constructed for the next predicted transaction. 
  typedef decode_out_transaction decode_out_ap_output_transaction_t;
  decode_out_ap_output_transaction_t decode_out_ap_output_transaction;
  // Code for sending output transaction out through decode_out_ap
  // decode_out_ap.write(decode_out_ap_output_transaction);

  // Define transaction handles for debug visibility 
  decode_in_transaction decode_in_ae_debug;


  // pragma uvmf custom class_item_additional begin
  // pragma uvmf custom class_item_additional end

  // FUNCTION: new
  function new(string name, uvm_component parent);
     super.new(name,parent);
    //`uvm_warning("PREDICTOR_REVIEW", "This predictor has been created either through generation or re-generation with merging.  Remove this warning after the predictor has been reviewed.")
  // pragma uvmf custom new begin
  // pragma uvmf custom new end
  endfunction

  // FUNCTION: build_phase
  virtual function void build_phase (uvm_phase phase);

    decode_in_ae = new("decode_in_ae", this);
    decode_out_ap =new("decode_out_ap", this );
  // pragma uvmf custom build_phase begin
  // pragma uvmf custom build_phase end
  endfunction

  // FUNCTION: write_decode_in_ae
  // Transactions received through decode_in_ae initiate the execution of this function.
  // This function performs prediction of DUT output values based on DUT input, configuration and state
  virtual function void write_decode_in_ae(decode_in_transaction t);
    // pragma uvmf custom decode_in_ae_predictor begin
    bit [15:0] ir, npc_out;
    bit [5:0] e_control;
    bit [1:0] w_control;
    bit mem_control;
    bit decode_model_output;

    //Harry: skip the prediction if the enable_decode is 0 since the actual output is not valid to compare with
    if (!t.enable_decode) begin
      `uvm_info("DECODE_PRED",
        $sformatf("Skipping decode prediction at %0t because enable_decode=0", $time),
        UVM_HIGH)
      return;
    end

    decode_in_ae_debug = t;
    

    /*decode_in_transaction
  rand bit [15:0] npc_in ;
  rand bit [15:0] instr_dout ;
  time start_time ;
  time end_time ;
  rand bit [3:0] psr ;
  rand bit enable_decode ;
    */
    `uvm_info("PRED", "Transaction Received through decode_in_ae", UVM_MEDIUM)
    `uvm_info("PRED", {"            Data: ",t.convert2string()}, UVM_FULL)
    // Construct one of each output transaction type.
    decode_out_ap_output_transaction = decode_out_ap_output_transaction_t::type_id::create("decode_out_ap_output_transaction");
    //  UVMF_CHANGE_ME: Implement predictor model here.  
    decode_model_output = decode_model(
      t.instr_dout, // input bit [15: 0] instr_dout,
      t.npc_in,     // input bit [15: 0] npc_in,
      ir,           // output bit [15: 0] ir,
      npc_out,      // output bit [15: 0] npc_out,
      e_control,    // output bit [5: 0] e_control,
      w_control,    // output bit [1: 0] w_control,
      mem_control   // output bit mem_control
    );

    decode_out_ap_output_transaction.ir = ir;
    decode_out_ap_output_transaction.npc_out = npc_out;
    decode_out_ap_output_transaction.e_control = e_control;
    decode_out_ap_output_transaction.w_control = w_control;
    decode_out_ap_output_transaction.mem_control = mem_control;

    // Code for sending output transaction out through decode_out_ap
    // Please note that each broadcasted transaction should be a different object than previously 
    // broadcasted transactions.  Creation of a different object is done by constructing the transaction 
    // using either new() or create().  Broadcasting a transaction object more than once to either the 
    // same subscriber or multiple subscribers will result in unexpected and incorrect behavior.
    decode_out_ap.write(decode_out_ap_output_transaction);
    `uvm_info("PRED", $sformatf("Prediction sent from decode_model: ir=0x%0h npc_out=0x%0h e_control=0x%0h w_control=0x%0h mem_control=0x%0h",
                            ir, npc_out, e_control, w_control, mem_control),
          UVM_LOW)
    // pragma uvmf custom decode_in_ae_predictor end
  endfunction

endclass

// pragma uvmf custom external begin
// pragma uvmf custom external end
