`define CPU_PC_COUNTER_SIZE 32
`define CPU_PC_NUMBER_OF_TRIGGERS 3
