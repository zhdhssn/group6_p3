//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4_2
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef bit [5:0] e_control_t;
typedef bit [15:0] ir_t;
typedef bit [15:0] npc_in_t;
typedef bit bypass_alu_1_t;
typedef bit bypass_alu_2_t;
typedef bit bypass_mem_1_t;
typedef bit bypass_mem_2_t;
typedef bit [15:0] vsr1_t;
typedef bit [15:0] vsr2_t;
typedef bit [1:0] w_control_in_t;
typedef bit mem_control_in_t;
typedef bit enable_execute_t;
typedef bit [15:0] mem_bypass_val_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

