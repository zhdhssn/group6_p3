package signal_monitor_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  //Include the components
  `include "signal_monitor_proxy.svh"

endpackage : signal_monitor_pkg


