package signal_driver_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  //Include the components
  `include "signal_driver_proxy.svh"

endpackage : signal_driver_pkg

