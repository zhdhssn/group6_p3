//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4_2
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: 
// This file contains defines and typedefs to be compiled for use in
// the simulation running on the emulator when using Veloce.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
                                                                               

typedef bit [1:0] w_control_out_t;
typedef bit mem_control_out_t;
typedef bit [15:0] aluout_t;
typedef bit [15:0] pcout_t;
typedef bit [2:0] dr_t;
typedef bit [2:0] sr1_t;
typedef bit [2:0] sr2_t;
typedef bit [15:0] ir_exec_t;
typedef bit [2:0] nzp_t;
typedef bit [15:0] m_data_t;
typedef bit enable_execute_t;

// pragma uvmf custom additional begin
// pragma uvmf custom additional end

